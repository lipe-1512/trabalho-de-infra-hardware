module mux_memory_reg (
    ports
);
    
endmodule