module moduleName (
    input wire clk, reset,
    input wire 0, OpCode, F
);
    
endmodule